module instMem(   //as rom memory
    input logic [10:0] i_addr,
    output logic [31:0] o_data
);
logic [7:0] mem [0: 2047]; //intermal memory block

assign mem[0] = 8'hb7;
assign mem[1] = 8'h3f;
assign mem[2] = 8'h00;
assign mem[3] = 8'h10;
assign mem[4] = 8'h37;
assign mem[5] = 8'h2f;
assign mem[6] = 8'h00;
assign mem[7] = 8'h10;
assign mem[8] = 8'hb7;
assign mem[9] = 8'h0e;
assign mem[10] = 8'h01;
assign mem[11] = 8'h10;
assign mem[12] = 8'h17;
assign mem[13] = 8'h0b;
assign mem[14] = 8'h00;
assign mem[15] = 8'h00;
assign mem[16] = 8'h13;
assign mem[17] = 8'h0b;
assign mem[18] = 8'hcb;
assign mem[19] = 8'h0d;
assign mem[20] = 8'h97;
assign mem[21] = 8'h0a;
assign mem[22] = 8'h00;
assign mem[23] = 8'h00;
assign mem[24] = 8'h93;
assign mem[25] = 8'h8a;
assign mem[26] = 8'h8a;
assign mem[27] = 8'h0b;
assign mem[28] = 8'hb7;
assign mem[29] = 8'h0d;
assign mem[30] = 8'h00;
assign mem[31] = 8'h10;
assign mem[32] = 8'h93;
assign mem[33] = 8'h0c;
assign mem[34] = 8'hf0;
assign mem[35] = 8'hff;
assign mem[36] = 8'hb7;
assign mem[37] = 8'hf1;
assign mem[38] = 8'hfa;
assign mem[39] = 8'h02;
assign mem[40] = 8'h93;
assign mem[41] = 8'h81;
assign mem[42] = 8'h01;
assign mem[43] = 8'h08;
assign mem[44] = 8'h13;
assign mem[45] = 8'h02;
assign mem[46] = 8'hc0;
assign mem[47] = 8'h03;
assign mem[48] = 8'h93;
assign mem[49] = 8'h00;
assign mem[50] = 8'h10;
assign mem[51] = 8'h00;
assign mem[52] = 8'h13;
assign mem[53] = 8'h01;
assign mem[54] = 8'h00;
assign mem[55] = 8'h00;
assign mem[56] = 8'h03;
assign mem[57] = 8'hae;
assign mem[58] = 8'h0e;
assign mem[59] = 8'h00;
assign mem[60] = 8'h13;
assign mem[61] = 8'h1e;
assign mem[62] = 8'h0e;
assign mem[63] = 8'h01;
assign mem[64] = 8'h13;
assign mem[65] = 8'h7e;
assign mem[66] = 8'h1e;
assign mem[67] = 8'h00;
assign mem[68] = 8'h63;
assign mem[69] = 8'h08;
assign mem[70] = 8'h0e;
assign mem[71] = 8'h00;
assign mem[72] = 8'h03;
assign mem[73] = 8'hae;
assign mem[74] = 8'h0e;
assign mem[75] = 8'h00;
assign mem[76] = 8'h93;
assign mem[77] = 8'h70;
assign mem[78] = 8'hfe;
assign mem[79] = 8'h00;
assign mem[80] = 8'h6f;
assign mem[81] = 8'hf0;
assign mem[82] = 8'h9f;
assign mem[83] = 8'hfe;
assign mem[84] = 8'h23;
assign mem[85] = 8'ha0;
assign mem[86] = 8'h0d;
assign mem[87] = 8'h00;
assign mem[88] = 8'h13;
assign mem[89] = 8'h85;
assign mem[90] = 8'h00;
assign mem[91] = 8'h00;
assign mem[92] = 8'h67;
assign mem[93] = 8'h8a;
assign mem[94] = 8'h0a;
assign mem[95] = 8'h00;
assign mem[96] = 8'h33;
assign mem[97] = 8'h8e;
assign mem[98] = 8'h65;
assign mem[99] = 8'h01;
assign mem[100] = 8'h03;
assign mem[101] = 8'h2e;
assign mem[102] = 8'h0e;
assign mem[103] = 8'h00;
assign mem[104] = 8'ha3;
assign mem[105] = 8'h80;
assign mem[106] = 8'hcf;
assign mem[107] = 8'h01;
assign mem[108] = 8'h33;
assign mem[109] = 8'h0e;
assign mem[110] = 8'h65;
assign mem[111] = 8'h01;
assign mem[112] = 8'h03;
assign mem[113] = 8'h2e;
assign mem[114] = 8'h0e;
assign mem[115] = 8'h00;
assign mem[116] = 8'h23;
assign mem[117] = 8'h80;
assign mem[118] = 8'hcf;
assign mem[119] = 8'h01;
assign mem[120] = 8'h13;
assign mem[121] = 8'h05;
assign mem[122] = 8'h01;
assign mem[123] = 8'h00;
assign mem[124] = 8'h67;
assign mem[125] = 8'h8a;
assign mem[126] = 8'h0a;
assign mem[127] = 8'h00;
assign mem[128] = 8'h33;
assign mem[129] = 8'h8e;
assign mem[130] = 8'h65;
assign mem[131] = 8'h01;
assign mem[132] = 8'h03;
assign mem[133] = 8'h2e;
assign mem[134] = 8'h0e;
assign mem[135] = 8'h00;
assign mem[136] = 8'ha3;
assign mem[137] = 8'h00;
assign mem[138] = 8'hcf;
assign mem[139] = 8'h01;
assign mem[140] = 8'h33;
assign mem[141] = 8'h0e;
assign mem[142] = 8'h65;
assign mem[143] = 8'h01;
assign mem[144] = 8'h03;
assign mem[145] = 8'h2e;
assign mem[146] = 8'h0e;
assign mem[147] = 8'h00;
assign mem[148] = 8'h23;
assign mem[149] = 8'h00;
assign mem[150] = 8'hcf;
assign mem[151] = 8'h01;
assign mem[152] = 8'h63;
assign mem[153] = 8'h0e;
assign mem[154] = 8'h01;
assign mem[155] = 8'h00;
assign mem[156] = 8'h63;
assign mem[157] = 8'h86;
assign mem[158] = 8'h32;
assign mem[159] = 8'h00;
assign mem[160] = 8'h93;
assign mem[161] = 8'h82;
assign mem[162] = 8'h12;
assign mem[163] = 8'h00;
assign mem[164] = 8'h6f;
assign mem[165] = 8'hf0;
assign mem[166] = 8'h9f;
assign mem[167] = 8'hff;
assign mem[168] = 8'h93;
assign mem[169] = 8'h02;
assign mem[170] = 8'h00;
assign mem[171] = 8'h00;
assign mem[172] = 8'h13;
assign mem[173] = 8'h01;
assign mem[174] = 8'hf1;
assign mem[175] = 8'hff;
assign mem[176] = 8'h6f;
assign mem[177] = 8'hf0;
assign mem[178] = 8'h5f;
assign mem[179] = 8'hfa;
assign mem[180] = 8'h63;
assign mem[181] = 8'h88;
assign mem[182] = 8'h00;
assign mem[183] = 8'h00;
assign mem[184] = 8'h93;
assign mem[185] = 8'h80;
assign mem[186] = 8'hf0;
assign mem[187] = 8'hff;
assign mem[188] = 8'h13;
assign mem[189] = 8'h01;
assign mem[190] = 8'hb0;
assign mem[191] = 8'h03;
assign mem[192] = 8'h6f;
assign mem[193] = 8'hf0;
assign mem[194] = 8'h5f;
assign mem[195] = 8'hf9;
assign mem[196] = 8'h23;
assign mem[197] = 8'ha0;
assign mem[198] = 8'h9d;
assign mem[199] = 8'h01;
assign mem[200] = 8'h6f;
assign mem[201] = 8'hf0;
assign mem[202] = 8'h1f;
assign mem[203] = 8'hf7;
assign mem[204] = 8'h93;
assign mem[205] = 8'h06;
assign mem[206] = 8'ha0;
assign mem[207] = 8'h00;
assign mem[208] = 8'h93;
assign mem[209] = 8'h05;
assign mem[210] = 8'h00;
assign mem[211] = 8'h00;
assign mem[212] = 8'h63;
assign mem[213] = 8'h54;
assign mem[214] = 8'hd5;
assign mem[215] = 8'h00;
assign mem[216] = 8'h67;
assign mem[217] = 8'h00;
assign mem[218] = 8'h0a;
assign mem[219] = 8'h00;
assign mem[220] = 8'h13;
assign mem[221] = 8'h05;
assign mem[222] = 8'h65;
assign mem[223] = 8'hff;
assign mem[224] = 8'h93;
assign mem[225] = 8'h85;
assign mem[226] = 8'h15;
assign mem[227] = 8'h00;
assign mem[228] = 8'h6f;
assign mem[229] = 8'hf0;
assign mem[230] = 8'h1f;
assign mem[231] = 8'hff;
assign mem[232] = 8'h40;
assign mem[233] = 8'h00;
assign mem[234] = 8'h00;
assign mem[235] = 8'h00;
assign mem[236] = 8'h79;
assign mem[237] = 8'h00;
assign mem[238] = 8'h00;
assign mem[239] = 8'h00;
assign mem[240] = 8'h24;
assign mem[241] = 8'h00;
assign mem[242] = 8'h00;
assign mem[243] = 8'h00;
assign mem[244] = 8'h30;
assign mem[245] = 8'h00;
assign mem[246] = 8'h00;
assign mem[247] = 8'h00;
assign mem[248] = 8'h19;
assign mem[249] = 8'h00;
assign mem[250] = 8'h00;
assign mem[251] = 8'h00;
assign mem[252] = 8'h12;
assign mem[253] = 8'h00;
assign mem[254] = 8'h00;
assign mem[255] = 8'h00;
assign mem[256] = 8'h02;
assign mem[257] = 8'h00;
assign mem[258] = 8'h00;
assign mem[259] = 8'h00;
assign mem[260] = 8'h78;
assign mem[261] = 8'h00;
assign mem[262] = 8'h00;
assign mem[263] = 8'h00;
assign mem[264] = 8'h00;
assign mem[265] = 8'h00;
assign mem[266] = 8'h00;
assign mem[267] = 8'h00;
assign mem[268] = 8'h10;
assign mem[269] = 8'h00;
assign mem[270] = 8'h00;
assign mem[271] = 8'h00;

logic [10:0] addr_0, addr_1, addr_2, addr_3;
assign addr_0 = i_addr;          // addr0 first byte
assign addr_1 = i_addr + 11'd1;  // addr1 second byte
assign addr_2 = i_addr + 11'd2;  // addr2 third byte
assign addr_3 = i_addr + 11'd3;  // addr3 four th byte
always @(*) begin
    o_data[7:0] = mem[addr_0];
    o_data[15:8] = mem[addr_1]; 
    o_data[23:16] = mem[addr_2];
    o_data[31:24] = mem[addr_3];  
end
endmodule